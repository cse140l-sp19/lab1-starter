//
// Lab1_hello
// CSE140L Spring 2019
//
// Starter code
//   Bryan Chin
//   Lih-Feng Tsaur
//
// Author:
//

module Lab1_hello(input tb_a, input tb_b, input tb_c, output L1_andOut);

   //Example boolean operation
   assign L1_andOut = tb_a & tb_b & tb_c;
   

endmodule

//
// Lab1_hello
// CSE140L Spring 2019
//
// Starter code
//   Bryan Chin
//   Lih-Feng Tsaur
//
// Author:
//

module Lab1_hello(input tb_a, input tb_b, output L1_c_a_and_b);

   assign L1_c_a_and_b = a & b;

endmodule

//
// Lab1_hello
// CSE140L Spring 2019
//
// Starter code
//   Bryan Chin
//   Lih-Feng Tsaur
//
// Author:
//

module Lab1_hello(input a, input b, output c_a_and_b);

   assign c_a_and_b = a & b;

endmodule
